

class test_zynq_class;
	

	
endclass : test_zynq_class
